`timescale 1 ns/1 ps

module fsm_mux_tb;

reg [13:0] U0 = 14'b00101001110110;
reg [13:0] U1 = 14'b00011101010100;
reg [13:0] U0_p = 14'b00000000000111;
reg [13:0] U0_m = 14'b11111111111001;
reg [13:0] U1_p = 14'b11111111111000;
reg [13:0] U1_m = 14'b00000000000101;

wire [13:0] DAC_A;
wire [13:0] DAC_B;

reg ADC_CLK;
wire [1:0] DAC_SEL;
reg TRIG_IN;
reg start = 1;

localparam ADC_CLK_HPERIOD = 2;
localparam TRIG_CLK_HPERIOD = 40;

DAC_MUX #(.DATA_WIDTH(14)) DAC_CON(.adc_clk(ADC_CLK), .DAC_SEL(DAC_SEL), .U0(U0), .U1(U1), .U0_p(U0_p), .U0_m(U0_m), .U1_p(U1_p), .U1_m(U1_m), .DAC_A_OUT(DAC_A), .DAC_B_OUT(DAC_B));

FSM CON_BOX(.TRIG_IN(TRIG_IN), .adc_clk(ADC_CLK), .start(start), .FSM_ADC_COUNTER_TRIG(FSM_ADC_COUNTER_TRIG), .FSM_DAC_COUNTER_TRIG(FSM_DAC_COUNTER_TRIG), .FSM_JP_WRT(), 
.FSM_JM_WRT(), .FSM_REG_RST(), .FSM_U_WRT(), .FSM_DAC_SEL(DAC_SEL), .FSM_ADC_COUNTER_START(FSM_ADC_COUNTER_START), .FSM_ADC_COUNTER_RST(FSM_ADC_COUNTER_RST),
.FSM_DAC_COUNTER_START(FSM_DAC_COUNTER_START), .FSM_DAC_COUNTER_RST(FSM_DAC_COUNTER_RST));

gen_counter #(.COUNT_DATA_WIDTH(4), .COUNTER_TRIG_VAL(10)) ADC_SAMP_COUNTER(.clk(ADC_CLK), .rst(FSM_ADC_COUNTER_RST), .en(FSM_ADC_COUNTER_START), .f(FSM_ADC_COUNTER_TRIG));
gen_counter #(.COUNT_DATA_WIDTH(4), .COUNTER_TRIG_VAL(7)) DAC_SAMP_COUNTER(.clk(ADC_CLK), .rst(FSM_DAC_COUNTER_RST), .en(FSM_DAC_COUNTER_START), .f(FSM_DAC_COUNTER_TRIG));

	always 
	begin
		ADC_CLK = 1'b0; 
		#ADC_CLK_HPERIOD;
		ADC_CLK = 1'b1;
		#ADC_CLK_HPERIOD;
	end
	always 
	begin
		TRIG_IN = 1'b0; 
		#TRIG_CLK_HPERIOD;
		TRIG_IN = 1'b1;
		#TRIG_CLK_HPERIOD;
	end

	initial
	begin
		#TRIG_CLK_HPERIOD;
		
	end
endmodule
