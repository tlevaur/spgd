module GPIO_PARAMS_WRAPPER #(
	parameter GPIO_WIDTH = 32,
	parameter PARAM_COUNT = 16,
	parameter PARAM_SETS = 16
)(
	input [PARAM_COUNT*(GPIO_WIDTH - 1)*PARAM_SETS: 0] PARAMS_DATA,
	input [3:0] SET,
	output [GPIO_WIDTH - 1 : 0] GP_OUT
);
	// GPIO Parameter Setup
	reg [GPIO_WIDTH - 1 : 0] GP_OUT_SET = {GPIO_WIDTH{1'b0}};
	assign GP_OUT = GP_OUT_SET; 

	localparam [3:0]
		GP_OUT_PARAM_SET0 = 4'h0,
		GP_OUT_PARAM_SET1 = 4'h1,
		GP_OUT_PARAM_SET2 = 4'h2,
		GP_OUT_PARAM_SET3 = 4'h3,
		GP_OUT_PARAM_SET4 = 4'h4,
		GP_OUT_PARAM_SET5 = 4'h5,
		GP_OUT_PARAM_SET6 = 4'h6,
		GP_OUT_PARAM_SET7 = 4'h7,
		GP_OUT_PARAM_SET8 = 4'h8,
		GP_OUT_PARAM_SET9 = 4'h9,
		GP_OUT_PARAM_SET10 = 4'hA,
		GP_OUT_PARAM_SET11 = 4'hB,
		GP_OUT_PARAM_SET12 = 4'hC,
		GP_OUT_PARAM_SET13 = 4'hD,
		GP_OUT_PARAM_SET14 = 4'hE,
		GP_OUT_PARAM_SET15 = 4'hF;

	always @(PARAMS_DATA or SET)
		begin
			case(SET)
				GP_OUT_PARAM_SET0 : GP_OUT_SET = PARAMS_DATA[PARAM_COUNT * GPIO_WIDTH *  1 - 1 : PARAM_COUNT * GPIO_WIDTH *  0];
				GP_OUT_PARAM_SET1 : GP_OUT_SET = PARAMS_DATA[PARAM_COUNT * GPIO_WIDTH *  2 - 1 : PARAM_COUNT * GPIO_WIDTH *  1];
				GP_OUT_PARAM_SET2 : GP_OUT_SET = PARAMS_DATA[PARAM_COUNT * GPIO_WIDTH *  3 - 1 : PARAM_COUNT * GPIO_WIDTH *  2];
				GP_OUT_PARAM_SET3 : GP_OUT_SET = PARAMS_DATA[PARAM_COUNT * GPIO_WIDTH *  4 - 1 : PARAM_COUNT * GPIO_WIDTH *  3];
				GP_OUT_PARAM_SET4 : GP_OUT_SET = PARAMS_DATA[PARAM_COUNT * GPIO_WIDTH *  5 - 1 : PARAM_COUNT * GPIO_WIDTH *  4];
				GP_OUT_PARAM_SET5 : GP_OUT_SET = PARAMS_DATA[PARAM_COUNT * GPIO_WIDTH *  6 - 1 : PARAM_COUNT * GPIO_WIDTH *  5];
				GP_OUT_PARAM_SET6 : GP_OUT_SET = PARAMS_DATA[PARAM_COUNT * GPIO_WIDTH *  7 - 1 : PARAM_COUNT * GPIO_WIDTH *  6];
				GP_OUT_PARAM_SET7 : GP_OUT_SET = PARAMS_DATA[PARAM_COUNT * GPIO_WIDTH *  8 - 1 : PARAM_COUNT * GPIO_WIDTH *  7];
				GP_OUT_PARAM_SET8 : GP_OUT_SET = PARAMS_DATA[PARAM_COUNT * GPIO_WIDTH *  9 - 1 : PARAM_COUNT * GPIO_WIDTH *  8];
				GP_OUT_PARAM_SET9 : GP_OUT_SET = PARAMS_DATA[PARAM_COUNT * GPIO_WIDTH * 10 - 1 : PARAM_COUNT * GPIO_WIDTH *  9];
				GP_OUT_PARAM_SET10: GP_OUT_SET = PARAMS_DATA[PARAM_COUNT * GPIO_WIDTH * 11 - 1 : PARAM_COUNT * GPIO_WIDTH * 10];
				GP_OUT_PARAM_SET11: GP_OUT_SET = PARAMS_DATA[PARAM_COUNT * GPIO_WIDTH * 12 - 1 : PARAM_COUNT * GPIO_WIDTH * 11];
				GP_OUT_PARAM_SET12: GP_OUT_SET = PARAMS_DATA[PARAM_COUNT * GPIO_WIDTH * 13 - 1 : PARAM_COUNT * GPIO_WIDTH * 12];
				GP_OUT_PARAM_SET13: GP_OUT_SET = PARAMS_DATA[PARAM_COUNT * GPIO_WIDTH * 14 - 1 : PARAM_COUNT * GPIO_WIDTH * 13];
				GP_OUT_PARAM_SET14: GP_OUT_SET = PARAMS_DATA[PARAM_COUNT * GPIO_WIDTH * 15 - 1 : PARAM_COUNT * GPIO_WIDTH * 14];
				GP_OUT_PARAM_SET15: GP_OUT_SET = PARAMS_DATA[PARAM_COUNT * GPIO_WIDTH * 16 - 1 : PARAM_COUNT * GPIO_WIDTH * 15];
				default		  : GP_OUT_SET = PARAMS_DATA[PARAM_COUNT * GPIO_WIDTH *  1 - 1 : PARAM_COUNT * GPIO_WIDTH *  0];
			endcase
		end
endmodule