module new_FSM_tb;

reg TRIG_IN = 1'b0;
reg adc_clk = 1'b0;
reg start = 1'b0;
wire FSM_JP_WRT;
wire FSM_JM_WRT;
wire FSM_U_WRT;
wire [1:0] FSM_DAC_SEL;
wire [5:0] FSM_STATE;


new_FSM FSM(.TRIG_IN(TRIG_IN), .adc_clk(adc_clk), .start(start), .FSM_JP_WRT(FSM_JP_WRT), .FSM_JM_WRT(FSM_JM_WRT), .FSM_U_WRT(FSM_U_WRT), .FSM_DAC_SEL(FSM_DAC_SEL), .FSM_STATE(FSM_STATE));

initial
begin
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	start = 1'b1;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	TRIG_IN = 1'b1;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	TRIG_IN = 1'b0;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 adc_clk = ~adc_clk;
	#10 $finish;
end
endmodule
