module CON_ORS
(
	input F_JP_WRT,
	input G_JP_WRT,
	input F_JM_WRT,
	input G_JP_WRT,
	input F_U_WRT,
	input G_U_WRT,
	output JP_WRT,
	output JM_WRT,
	output U_WRT,
)

endmodule
